`include "defines.v"

module ex_mem(

);

endmodule
