`include "defines.h"

module div(

);

endmodule
