`include "defines.v"

module mem_wb(

);

endmodule
