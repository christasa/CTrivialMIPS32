`include "defines.v"

module mem(


);

endmodule
