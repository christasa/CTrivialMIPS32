`include "defines.v"

module ex(

);

endmodule
