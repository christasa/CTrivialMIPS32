`include "defines.v"

module if_id(

);

endmodule