`include "defines.v"

module id_ex(

);

endmodule